module control_unit(
	input [5:0] opcode,
	input [5:0] funct,
	output reg [3:0] ALU_Code,
	output reg [1:0] regDst,
	output reg regWrite,
   output reg branch,
   output reg condZero,
   output reg aluSrc,
	output reg memWrite,
   output reg [1:0] memToReg,
   output reg [1:0] pcSrc
);	
always @(*) begin
	if (opcode == 6'b001001 || opcode == 6'b001100 || opcode == 6'b001101 || opcode == 6'b001011 || opcode == 6'b001111) begin
		regDst = 2'b00;
		regWrite = 1;
		branch = 0;
		condZero = 0;
		aluSrc = 1;
		memWrite = 0;
		memToReg = 2'b00;
		pcSrc = 2'b00;
		case (opcode)
			6'b001001: ALU_Code = 4'b0101;
			6'b001100: ALU_Code = 4'b0001;
			6'b001101: ALU_Code = 4'b0011;
			6'b001011: ALU_Code = 4'b1000;
			6'b001111: ALU_Code = 4'b1100;
		endcase
	end
	case (opcode)
		6'b000000: begin 
			regDst = 2'b01;
			regWrite = 1;
			branch = 0;
			condZero = 0;
			aluSrc = 0;
			memWrite = 0;
			memToReg = 2'b00;
			pcSrc = 2'b00;
			case (funct)
				6'b100001: ALU_Code = 4'b0101;
				6'b100011: ALU_Code = 4'b0110;
				6'b100100: ALU_Code = 4'b0001;
				6'b100101: ALU_Code = 4'b0011;
				6'b100110: ALU_Code = 4'b0010;
				6'b101011: ALU_Code = 4'b1000;
				6'b000000: ALU_Code = 4'b1010;
				6'b000010: ALU_Code = 4'b1010;
				6'b001000: begin 
					ALU_Code = 4'b0110;
					regWrite = 0;
					pcSrc = 2'b10;
				end
			endcase
		end
		6'b000100: begin
			ALU_Code = 4'b0110;
			regDst = 2'b00;
			regWrite = 0;
			branch = 1;
			condZero = 1;
			aluSrc = 1;
			memWrite = 0;
			memToReg = 2'b00;
			pcSrc = 2'b00;
		end
		6'b000101: begin
			ALU_Code = 4'b0110;
			regDst = 2'b00;
			regWrite = 0;
			branch = 1;
			condZero = 0;
			aluSrc = 1;
			memWrite = 0;
			memToReg = 2'b00;
			pcSrc = 2'b00;
		end
		6'b100011: begin
			ALU_Code = 4'b0101;
			regDst = 2'b00;
			regWrite = 1;
			branch = 0;
			condZero = 0;
			aluSrc = 1;
			memWrite = 0;
			memToReg = 2'b01;
			pcSrc = 2'b00;
		end
		6'b101011: begin
			ALU_Code = 4'b0101;
			regDst = 2'b00;
			regWrite = 0;
			branch = 0;
			condZero = 0;
			aluSrc = 1;
			memWrite = 1;
			memToReg = 2'b00;
			pcSrc = 2'b00;
		end
		6'b000010: begin
			ALU_Code = 4'b0110;
			regDst = 2'b00;
			regWrite = 0;
			branch = 0;
			condZero = 0;
			aluSrc = 0;
			memWrite = 0;
			memToReg = 2'b00;
			pcSrc = 2'b01;
		end
		6'b000011: begin
			ALU_Code = 4'b0110;
			regDst = 2'b10;
			regWrite = 1;
			branch = 0;
			condZero = 0;
			aluSrc = 0;
			memWrite = 0;
			memToReg = 2'b10;
			pcSrc = 2'b01;
		end
	endcase
end
endmodule
		
			
				